001
00b
800
111
113
800
011
013
800
081
083
000
181
183
800
