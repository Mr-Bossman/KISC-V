01
03
0b
00
11
13
00
