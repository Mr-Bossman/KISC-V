001
003
00b
000
011
013
000
081
083
181
183
000
