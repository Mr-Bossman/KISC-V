010001
02000b
000000
000000
000000
000000
000000
000000
090010
0a0015
0b0017
000000
000000
000000
000000
000000
110010
120011
130013
000000
000000
000000
000000
000000
190080
1a0081
1b0083
1c0000
1d0085
1e0087
000000
000000
210100
000000
000000
000000
000000
000000
000000
000000
290040
000000
000000
000000
000000
000000
000000
000000
310020
000000
000000
000000
000000
000000
000000
000000
000200
000000
000000
000000
000000
000000
000000
000000
000400
000000
000000
000000
000000
000000
000000
000000
