01
03
0b
00
04
00
00
00
11
13
00
00
00
