000001
00000b
000800
000000
000000
000000
000000
000000
000010
000111
000113
000800
000000
000000
000000
000000
000010
000011
000013
000800
000000
000000
000000
000000
000081
000083
000000
000181
000183
000800
000000
000000
000004
000800
000000
000000
000000
000000
000000
000000
000040
000800
000000
000000
000000
000000
000000
000000
000020
000800
000000
000000
000000
000000
000000
000000
000800
000000
000000
000000
000000
000000
000000
000000
000800
000000
000000
000000
000000
000000
000000
000000
